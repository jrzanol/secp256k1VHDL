LIBRARY ieee;
USE ieee.std_logic_1164.all;

PACKAGE MYWORK IS

CONSTANT P : STD_LOGIC_VECTOR (255 DOWNTO 0) := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFC2F";
CONSTANT Gx : STD_LOGIC_VECTOR (255 DOWNTO 0) := X"79BE667EF9DCBBAC55A06295CE870B07029BFCDB2DCE28D959F2815B16F81798";
CONSTANT Gy : STD_LOGIC_VECTOR (255 DOWNTO 0) := X"483ADA7726A3C4655DA4FBFC0E1108A8FD17B448A68554199C47D08FFB10D4B8";

COMPONENT secp256k1_AddOnePoint IS
PORT(Clock, Reset: IN STD_LOGIC;
		X1, Y1: IN STD_LOGIC_VECTOR (255 DOWNTO 0);
		XOUT, YOUT: OUT STD_LOGIC_VECTOR (255 DOWNTO 0);
		SignalOut: OUT STD_LOGIC);
END COMPONENT;

COMPONENT secp256k1_ModAdd IS
PORT(X1, X2: IN STD_LOGIC_VECTOR (255 DOWNTO 0);
		XOUT: OUT STD_LOGIC_VECTOR (255 DOWNTO 0));
END COMPONENT;

COMPONENT secp256k1_ModSub IS
PORT(X1, X2: IN STD_LOGIC_VECTOR (255 DOWNTO 0);
		XOUT: OUT STD_LOGIC_VECTOR (255 DOWNTO 0));
END COMPONENT;

COMPONENT secp256k1_ModMult IS
PORT(A, B: IN STD_LOGIC_VECTOR(255 DOWNTO 0);
		XOUT: OUT STD_LOGIC_VECTOR(255 DOWNTO 0));
END COMPONENT;

COMPONENT secp256k1_ModNeg IS
PORT(X1: IN STD_LOGIC_VECTOR (255 DOWNTO 0);
		XOUT: OUT STD_LOGIC_VECTOR (255 DOWNTO 0));
END COMPONENT;

END PACKAGE;

